module regfile(
    input         clk,
    // READ PORT 1
    input  [ 4:0] raddr1,//共32个64位寄存器
    output [63:0] rdata1,
    // READ PORT 2
    input  [ 4:0] raddr2,
    output [63:0] rdata2,
    // WRITE PORT
    input         we,       //
    input  [ 4:0] waddr,
    input  [63:0] wdata

    // output [63:0] debug_rdata1,
    // output [63:0] debug_rdata2,
);
reg [63:0] rf[31:0];


always @(posedge clk) begin
    if (we) rf[waddr]<= wdata;
end


assign rdata1 = (raddr1==5'b0) ? 64'b0 : rf[raddr1];

assign rdata2 = (raddr2==5'b0) ? 64'b0 : rf[raddr2];

// assign debug_rdata1 =rdata1;
// assign debug_rdata2 =rdata2;
endmodule